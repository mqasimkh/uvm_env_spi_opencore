class wish_sequence extends uvm_sequence#(wish_packet);
    `uvm_object_utils(wish_sequence)

    function new (string name = "wish_sequence");
        super.new(name);
    endfunction: new

    function void build_phase (uvm_phase phase);
        `uvm_info(get_type_name(), "BUILD PHASE RUNNING ...", UVM_LOW)
    endfunction: build_phase

  task pre_body();
    uvm_phase phase;
    `ifdef UVM_VERSION_1_2
      phase = get_starting_phase();
    `else
      phase = starting_phase;
    `endif
    if (phase != null) begin
      phase.raise_objection(this, get_type_name());
      `uvm_info(get_type_name(), "OBJECTION RAISED", UVM_MEDIUM)
    end
  endtask : pre_body

  task post_body();
    uvm_phase phase;
    `ifdef UVM_VERSION_1_2
      phase = get_starting_phase();
    `else
      phase = starting_phase;
    `endif
    if (phase != null) begin
      
      phase.drop_objection(this, get_type_name());
      `uvm_info(get_type_name(), "OBJECTION DROPPED", UVM_MEDIUM)
    end
  endtask : post_body

endclass: wish_sequence

////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////                         test_sequence                                      //////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

class test_sequence extends wish_sequence;
    `uvm_object_utils(test_sequence)

    function new (string name = "test_sequence");
        super.new(name);
    endfunction: new

    virtual task body();
        `uvm_info(get_type_name(), "Running Sequence test_sequence ...", UVM_LOW)
        repeat(5) begin
            `uvm_do(req)
        end
    endtask: body

endclass: test_sequence