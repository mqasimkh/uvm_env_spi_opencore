package wish_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "wish_packet.sv"

endpackage: wish_pkg