interface spis_if();

  logic sck_o,
  logic ss_o,
  logic mosi_o,
  logic miso_i    

endinterface: spis_if